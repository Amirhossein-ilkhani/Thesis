module Generator_Addr_in #(
	parameter ROW = 4,
	parameter COL = 4,
	ROW 
	)(
	input clk,rst,en,
	input [7:0] i,j,k,
	

	);
	

endmodule